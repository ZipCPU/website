
	// Taken from a much larger module
	input	wire	A;
	output	wire	B;

	OBUF obuf(.I(B), .O(A));




